// A simple AND function

module simpleand(f,x,y);

  input x,y;
  output f;
  assign f= x& y;

endmodule